library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package cpu_types is


  subtype rst_system is std_logic;
  type array_of_signed_12 is array (integer range <>) of signed(11 downto 0);
  type tup3 is record
    tup3_sel0_signed : signed(11 downto 0);
    tup3_sel1_array_of_signed_12_0 : cpu_types.array_of_signed_12(0 to 1);
    tup3_sel2_array_of_signed_12_1 : cpu_types.array_of_signed_12(0 to 15);
  end record;
  subtype clk_system is std_logic;
  function toSLV (b : in boolean) return std_logic_vector;
  function fromSLV (sl : in std_logic_vector) return boolean;
  function tagToEnum (s : in signed) return boolean;
  function dataToTag (b : in boolean) return signed;
  function toSLV (s : in signed) return std_logic_vector;
  function fromSLV (slv : in std_logic_vector) return signed;
  function toSLV (sl : in std_logic) return std_logic_vector;
  function fromSLV (slv : in std_logic_vector) return std_logic;
  function toSLV (value :  cpu_types.array_of_signed_12) return std_logic_vector;
  function fromSLV (slv : in std_logic_vector) return cpu_types.array_of_signed_12;
  function toSLV (p : cpu_types.tup3) return std_logic_vector;
  function fromSLV (slv : in std_logic_vector) return cpu_types.tup3;
end;

package body cpu_types is
  function toSLV (b : in boolean) return std_logic_vector is
  begin
    if b then
      return "1";
    else
      return "0";
    end if;
  end;
  function fromSLV (sl : in std_logic_vector) return boolean is
  begin
    if sl = "1" then
      return true;
    else
      return false;
    end if;
  end;
  function tagToEnum (s : in signed) return boolean is
  begin
    if s = to_signed(0,64) then
      return false;
    else
      return true;
    end if;
  end;
  function dataToTag (b : in boolean) return signed is
  begin
    if b then
      return to_signed(1,64);
    else
      return to_signed(0,64);
    end if;
  end;
  function toSLV (s : in signed) return std_logic_vector is
  begin
    return std_logic_vector(s);
  end;
  function fromSLV (slv : in std_logic_vector) return signed is
  begin
    return signed(slv);
  end;
  function toSLV (sl : in std_logic) return std_logic_vector is
  begin
    return std_logic_vector'(0 => sl);
  end;
  function fromSLV (slv : in std_logic_vector) return std_logic is
    alias islv : std_logic_vector (0 to slv'length - 1) is slv;
  begin
    return islv(0);
  end;
  function toSLV (value :  cpu_types.array_of_signed_12) return std_logic_vector is
    alias ivalue    : cpu_types.array_of_signed_12(1 to value'length) is value;
    variable result : std_logic_vector(1 to value'length * 12);
  begin
    for i in ivalue'range loop
      result(((i - 1) * 12) + 1 to i*12) := toSLV(ivalue(i));
    end loop;
    return result;
  end;
  function fromSLV (slv : in std_logic_vector) return cpu_types.array_of_signed_12 is
    alias islv      : std_logic_vector(0 to slv'length - 1) is slv;
    variable result : cpu_types.array_of_signed_12(0 to slv'length / 12 - 1);
  begin
    for i in result'range loop
      result(i) := fromSLV(islv(i * 12 to (i+1) * 12 - 1));
    end loop;
    return result;
  end;
  function toSLV (p : cpu_types.tup3) return std_logic_vector is
  begin
    return (toSLV(p.tup3_sel0_signed) & toSLV(p.tup3_sel1_array_of_signed_12_0) & toSLV(p.tup3_sel2_array_of_signed_12_1));
  end;
  function fromSLV (slv : in std_logic_vector) return cpu_types.tup3 is
  alias islv : std_logic_vector(0 to slv'length - 1) is slv;
  begin
    return (fromSLV(islv(0 to 11)),fromSLV(islv(12 to 35)),fromSLV(islv(36 to 227)));
  end;
end;

